module Encoder_16x4(output reg [3:0] z, input [15:0] a);

always@(a)
begin
case(a)
16'b0000000000000001 : z  = 4'b0000;
16'b0000000000000010 : z  = 4'b0001;
16'b0000000000000100 : z  = 4'b0010;
16'b0000000000001000 : z  = 4'b0011;
16'b0000000000010000 : z  = 4'b0100;
16'b0000000000100000 : z  = 4'b0101;
16'b0000000001000000 : z  = 4'b0110;
16'b0000000010000000 : z  = 4'b0111;
16'b0000000100000000 : z  = 4'b1000;
16'b0000001000000000 : z  = 4'b1001;
16'b0000010000000000 : z  = 4'b1010;
16'b0000100000000000 : z  = 4'b1011;
16'b0001000000000000 : z  = 4'b1100;
16'b0010000000000000 : z  = 4'b1101;
16'b0100000000000000 : z  = 4'b1110;
16'b1000000000000000 : z  = 4'b1111;

default : z = 4'bxxxx;
endcase
end
endmodule 

module Encoder_16x4_tb();
reg [15:0] a;
wire [3:0] z;

Encoder_16x4 DUT(z,a);

initial
begin

a = 16'b0000000000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000000000001; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000000000010; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000000000100; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000000001000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000000010000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000000100000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000001000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000010000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000000100000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000001000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000010000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0000100000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0001000000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0010000000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b0100000000000000; #10;
$display ("z = %b, a = %b",z,a);

a = 16'b1000000000000000; #10;
$display ("z = %b, a = %b",z,a);

#20; $finish;
end
endmodule